-------------------------------------------------
-- File:	MUX.vhd
-- Entity:	Multiplexer for ALU
-- Architecture:	Structural
-- Author: John Judge
-- Created: 3/15/16
-- Modified: 3/15/16
-- VHDL'93
-- Description: The following is the entity and
--	behavioral description of a 16-bit variable shifter
-------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;



entity MUX is
end MUX;

architecture Behavioral of MUX is

begin


end Behavioral;

